module sid_coeffs
  (
	input             clk,
	input [10:0]      addr,
   output reg [15:0] val
  );

   reg [15:0]        coeff [0:2047];

   initial
     begin
		  coeff[0] <= 16'h02d5;
        coeff[1] <= 16'h02d5;
        coeff[2] <= 16'h02d5;
        coeff[3] <= 16'h02d5;
        coeff[4] <= 16'h02d5;
        coeff[5] <= 16'h02d5;
        coeff[6] <= 16'h02d5;
        coeff[7] <= 16'h02d5;
        coeff[8] <= 16'h02d5;
        coeff[9] <= 16'h02d5;
        coeff[10] <= 16'h02d5;
        coeff[11] <= 16'h02d5;
        coeff[12] <= 16'h02d5;
        coeff[13] <= 16'h02d5;
        coeff[14] <= 16'h02d5;
        coeff[15] <= 16'h02d5;
		  coeff[16] <= 16'h02d5;
        coeff[17] <= 16'h02d8;
        coeff[18] <= 16'h02d8;
        coeff[19] <= 16'h02d8;
        coeff[20] <= 16'h02d8;
        coeff[21] <= 16'h02d8;
        coeff[22] <= 16'h02d8;
        coeff[23] <= 16'h02d8;
        coeff[24] <= 16'h02d8;
        coeff[25] <= 16'h02d8;
        coeff[26] <= 16'h02d8;
        coeff[27] <= 16'h02d8;
        coeff[28] <= 16'h02d8;
        coeff[29] <= 16'h02d8;
        coeff[30] <= 16'h02d8;
        coeff[31] <= 16'h02d8;
        coeff[32] <= 16'h02d8;
        coeff[33] <= 16'h02d8;
        coeff[34] <= 16'h02db;
        coeff[35] <= 16'h02db;
        coeff[36] <= 16'h02db;
        coeff[37] <= 16'h02db;
        coeff[38] <= 16'h02db;
        coeff[39] <= 16'h02db;
        coeff[40] <= 16'h02db;
        coeff[41] <= 16'h02db;
        coeff[42] <= 16'h02db;
        coeff[43] <= 16'h02db;
        coeff[44] <= 16'h02db;
        coeff[45] <= 16'h02db;
        coeff[46] <= 16'h02db;
        coeff[47] <= 16'h02db;
        coeff[48] <= 16'h02db;
        coeff[49] <= 16'h02df;
        coeff[50] <= 16'h02df;
        coeff[51] <= 16'h02df;
        coeff[52] <= 16'h02df;
        coeff[53] <= 16'h02df;
        coeff[54] <= 16'h02df;
        coeff[55] <= 16'h02df;
        coeff[56] <= 16'h02df;
        coeff[57] <= 16'h02df;
        coeff[58] <= 16'h02df;
        coeff[59] <= 16'h02df;
        coeff[60] <= 16'h02df;
        coeff[61] <= 16'h02df;
        coeff[62] <= 16'h02df;
        coeff[63] <= 16'h02df;
        coeff[64] <= 16'h02e2;
        coeff[65] <= 16'h02e2;
        coeff[66] <= 16'h02e2;
        coeff[67] <= 16'h02e2;
        coeff[68] <= 16'h02e2;
        coeff[69] <= 16'h02e2;
        coeff[70] <= 16'h02e2;
        coeff[71] <= 16'h02e2;
        coeff[72] <= 16'h02e2;
        coeff[73] <= 16'h02e2;
        coeff[74] <= 16'h02e2;
        coeff[75] <= 16'h02e2;
        coeff[76] <= 16'h02e2;
        coeff[77] <= 16'h02e5;
        coeff[78] <= 16'h02e5;
        coeff[79] <= 16'h02e5;
        coeff[80] <= 16'h02e5;
        coeff[81] <= 16'h02e5;
        coeff[82] <= 16'h02e5;
        coeff[83] <= 16'h02e5;
        coeff[84] <= 16'h02e5;
        coeff[85] <= 16'h02e5;
        coeff[86] <= 16'h02e5;
        coeff[87] <= 16'h02e5;
        coeff[88] <= 16'h02e5;
        coeff[89] <= 16'h02e8;
        coeff[90] <= 16'h02e8;
        coeff[91] <= 16'h02e8;
        coeff[92] <= 16'h02e8;
        coeff[93] <= 16'h02e8;
        coeff[94] <= 16'h02e8;
        coeff[95] <= 16'h02e8;
        coeff[96] <= 16'h02e8;
        coeff[97] <= 16'h02e8;
        coeff[98] <= 16'h02e8;
        coeff[99] <= 16'h02e8;
        coeff[100] <= 16'h02ec;
        coeff[101] <= 16'h02ec;
        coeff[102] <= 16'h02ec;
        coeff[103] <= 16'h02ec;
        coeff[104] <= 16'h02ec;
        coeff[105] <= 16'h02ec;
        coeff[106] <= 16'h02ec;
        coeff[107] <= 16'h02ec;
        coeff[108] <= 16'h02ec;
        coeff[109] <= 16'h02ec;
        coeff[110] <= 16'h02ef;
        coeff[111] <= 16'h02ef;
        coeff[112] <= 16'h02ef;
        coeff[113] <= 16'h02ef;
        coeff[114] <= 16'h02ef;
        coeff[115] <= 16'h02ef;
        coeff[116] <= 16'h02ef;
        coeff[117] <= 16'h02ef;
        coeff[118] <= 16'h02ef;
        coeff[119] <= 16'h02ef;
        coeff[120] <= 16'h02f2;
        coeff[121] <= 16'h02f2;
        coeff[122] <= 16'h02f2;
        coeff[123] <= 16'h02f2;
        coeff[124] <= 16'h02f2;
        coeff[125] <= 16'h02f2;
        coeff[126] <= 16'h02f2;
        coeff[127] <= 16'h02f2;
        coeff[128] <= 16'h02f6;
        coeff[129] <= 16'h02f6;
        coeff[130] <= 16'h02f6;
        coeff[131] <= 16'h02f6;
        coeff[132] <= 16'h02f6;
        coeff[133] <= 16'h02f6;
        coeff[134] <= 16'h02f6;
        coeff[135] <= 16'h02f6;
        coeff[136] <= 16'h02f6;
        coeff[137] <= 16'h02f9;
        coeff[138] <= 16'h02f9;
        coeff[139] <= 16'h02f9;
        coeff[140] <= 16'h02f9;
        coeff[141] <= 16'h02f9;
        coeff[142] <= 16'h02f9;
        coeff[143] <= 16'h02f9;
        coeff[144] <= 16'h02f9;
        coeff[145] <= 16'h02f9;
        coeff[146] <= 16'h02fc;
        coeff[147] <= 16'h02fc;
        coeff[148] <= 16'h02fc;
        coeff[149] <= 16'h02fc;
        coeff[150] <= 16'h02fc;
        coeff[151] <= 16'h02fc;
        coeff[152] <= 16'h02fc;
        coeff[153] <= 16'h02fc;
        coeff[154] <= 16'h02fc;
        coeff[155] <= 16'h0300;
        coeff[156] <= 16'h0300;
        coeff[157] <= 16'h0300;
        coeff[158] <= 16'h0300;
        coeff[159] <= 16'h0300;
        coeff[160] <= 16'h0300;
        coeff[161] <= 16'h0300;
        coeff[162] <= 16'h0300;
        coeff[163] <= 16'h0300;
        coeff[164] <= 16'h0303;
        coeff[165] <= 16'h0303;
        coeff[166] <= 16'h0303;
        coeff[167] <= 16'h0303;
        coeff[168] <= 16'h0303;
        coeff[169] <= 16'h0303;
        coeff[170] <= 16'h0303;
        coeff[171] <= 16'h0303;
        coeff[172] <= 16'h0303;
        coeff[173] <= 16'h0306;
        coeff[174] <= 16'h0306;
        coeff[175] <= 16'h0306;
        coeff[176] <= 16'h0306;
        coeff[177] <= 16'h0306;
        coeff[178] <= 16'h0306;
        coeff[179] <= 16'h0306;
        coeff[180] <= 16'h0306;
        coeff[181] <= 16'h0309;
        coeff[182] <= 16'h0309;
        coeff[183] <= 16'h0309;
        coeff[184] <= 16'h0309;
        coeff[185] <= 16'h0309;
        coeff[186] <= 16'h0309;
        coeff[187] <= 16'h0309;
        coeff[188] <= 16'h0309;
        coeff[189] <= 16'h030d;
        coeff[190] <= 16'h030d;
        coeff[191] <= 16'h030d;
        coeff[192] <= 16'h030d;
        coeff[193] <= 16'h030d;
        coeff[194] <= 16'h030d;
        coeff[195] <= 16'h030d;
        coeff[196] <= 16'h0310;
        coeff[197] <= 16'h0310;
        coeff[198] <= 16'h0310;
        coeff[199] <= 16'h0310;
        coeff[200] <= 16'h0310;
        coeff[201] <= 16'h0310;
        coeff[202] <= 16'h0310;
        coeff[203] <= 16'h0313;
        coeff[204] <= 16'h0313;
        coeff[205] <= 16'h0313;
        coeff[206] <= 16'h0313;
        coeff[207] <= 16'h0313;
        coeff[208] <= 16'h0313;
        coeff[209] <= 16'h0317;
        coeff[210] <= 16'h0317;
        coeff[211] <= 16'h0317;
        coeff[212] <= 16'h0317;
        coeff[213] <= 16'h0317;
        coeff[214] <= 16'h0317;
        coeff[215] <= 16'h031a;
        coeff[216] <= 16'h031a;
        coeff[217] <= 16'h031a;
        coeff[218] <= 16'h031a;
        coeff[219] <= 16'h031a;
        coeff[220] <= 16'h031a;
        coeff[221] <= 16'h031d;
        coeff[222] <= 16'h031d;
        coeff[223] <= 16'h031d;
        coeff[224] <= 16'h031d;
        coeff[225] <= 16'h031d;
        coeff[226] <= 16'h0320;
        coeff[227] <= 16'h0320;
        coeff[228] <= 16'h0320;
        coeff[229] <= 16'h0320;
        coeff[230] <= 16'h0320;
        coeff[231] <= 16'h0324;
        coeff[232] <= 16'h0324;
        coeff[233] <= 16'h0324;
        coeff[234] <= 16'h0324;
        coeff[235] <= 16'h0324;
        coeff[236] <= 16'h0327;
        coeff[237] <= 16'h0327;
        coeff[238] <= 16'h0327;
        coeff[239] <= 16'h0327;
        coeff[240] <= 16'h0327;
        coeff[241] <= 16'h032a;
        coeff[242] <= 16'h032a;
        coeff[243] <= 16'h032a;
        coeff[244] <= 16'h032a;
        coeff[245] <= 16'h032e;
        coeff[246] <= 16'h032e;
        coeff[247] <= 16'h032e;
        coeff[248] <= 16'h032e;
        coeff[249] <= 16'h0331;
        coeff[250] <= 16'h0331;
        coeff[251] <= 16'h0331;
        coeff[252] <= 16'h0331;
        coeff[253] <= 16'h0334;
        coeff[254] <= 16'h0334;
        coeff[255] <= 16'h0334;
        coeff[256] <= 16'h0338;
        coeff[257] <= 16'h0338;
        coeff[258] <= 16'h0338;
        coeff[259] <= 16'h0338;
        coeff[260] <= 16'h033b;
        coeff[261] <= 16'h033b;
        coeff[262] <= 16'h033b;
        coeff[263] <= 16'h033b;
        coeff[264] <= 16'h033e;
        coeff[265] <= 16'h033e;
        coeff[266] <= 16'h033e;
        coeff[267] <= 16'h033e;
        coeff[268] <= 16'h0341;
        coeff[269] <= 16'h0341;
        coeff[270] <= 16'h0341;
        coeff[271] <= 16'h0345;
        coeff[272] <= 16'h0345;
        coeff[273] <= 16'h0345;
        coeff[274] <= 16'h0345;
        coeff[275] <= 16'h0348;
        coeff[276] <= 16'h0348;
        coeff[277] <= 16'h0348;
        coeff[278] <= 16'h0348;
        coeff[279] <= 16'h034b;
        coeff[280] <= 16'h034b;
        coeff[281] <= 16'h034b;
        coeff[282] <= 16'h034f;
        coeff[283] <= 16'h034f;
        coeff[284] <= 16'h034f;
        coeff[285] <= 16'h034f;
        coeff[286] <= 16'h0352;
        coeff[287] <= 16'h0352;
        coeff[288] <= 16'h0352;
        coeff[289] <= 16'h0355;
        coeff[290] <= 16'h0355;
        coeff[291] <= 16'h0355;
        coeff[292] <= 16'h0355;
        coeff[293] <= 16'h0358;
        coeff[294] <= 16'h0358;
        coeff[295] <= 16'h0358;
        coeff[296] <= 16'h035c;
        coeff[297] <= 16'h035c;
        coeff[298] <= 16'h035c;
        coeff[299] <= 16'h035c;
        coeff[300] <= 16'h035f;
        coeff[301] <= 16'h035f;
        coeff[302] <= 16'h035f;
        coeff[303] <= 16'h0362;
        coeff[304] <= 16'h0362;
        coeff[305] <= 16'h0362;
        coeff[306] <= 16'h0366;
        coeff[307] <= 16'h0366;
        coeff[308] <= 16'h0366;
        coeff[309] <= 16'h0369;
        coeff[310] <= 16'h0369;
        coeff[311] <= 16'h0369;
        coeff[312] <= 16'h036c;
        coeff[313] <= 16'h036c;
        coeff[314] <= 16'h036c;
        coeff[315] <= 16'h0370;
        coeff[316] <= 16'h0370;
        coeff[317] <= 16'h0370;
        coeff[318] <= 16'h0373;
        coeff[319] <= 16'h0373;
        coeff[320] <= 16'h0373;
        coeff[321] <= 16'h0376;
        coeff[322] <= 16'h0376;
        coeff[323] <= 16'h0376;
        coeff[324] <= 16'h0379;
        coeff[325] <= 16'h0379;
        coeff[326] <= 16'h0379;
        coeff[327] <= 16'h037d;
        coeff[328] <= 16'h037d;
        coeff[329] <= 16'h0380;
        coeff[330] <= 16'h0380;
        coeff[331] <= 16'h0380;
        coeff[332] <= 16'h0383;
        coeff[333] <= 16'h0383;
        coeff[334] <= 16'h0383;
        coeff[335] <= 16'h0387;
        coeff[336] <= 16'h0387;
        coeff[337] <= 16'h038a;
        coeff[338] <= 16'h038a;
        coeff[339] <= 16'h038d;
        coeff[340] <= 16'h038d;
        coeff[341] <= 16'h038d;
        coeff[342] <= 16'h0390;
        coeff[343] <= 16'h0390;
        coeff[344] <= 16'h0394;
        coeff[345] <= 16'h0394;
        coeff[346] <= 16'h0397;
        coeff[347] <= 16'h0397;
        coeff[348] <= 16'h0397;
        coeff[349] <= 16'h039a;
        coeff[350] <= 16'h039a;
        coeff[351] <= 16'h039e;
        coeff[352] <= 16'h039e;
        coeff[353] <= 16'h03a1;
        coeff[354] <= 16'h03a1;
        coeff[355] <= 16'h03a4;
        coeff[356] <= 16'h03a4;
        coeff[357] <= 16'h03a8;
        coeff[358] <= 16'h03a8;
        coeff[359] <= 16'h03ab;
        coeff[360] <= 16'h03ab;
        coeff[361] <= 16'h03ae;
        coeff[362] <= 16'h03ae;
        coeff[363] <= 16'h03b1;
        coeff[364] <= 16'h03b1;
        coeff[365] <= 16'h03b5;
        coeff[366] <= 16'h03b8;
        coeff[367] <= 16'h03b8;
        coeff[368] <= 16'h03bb;
        coeff[369] <= 16'h03bb;
        coeff[370] <= 16'h03bf;
        coeff[371] <= 16'h03bf;
        coeff[372] <= 16'h03c2;
        coeff[373] <= 16'h03c5;
        coeff[374] <= 16'h03c5;
        coeff[375] <= 16'h03c8;
        coeff[376] <= 16'h03c8;
        coeff[377] <= 16'h03cc;
        coeff[378] <= 16'h03cf;
        coeff[379] <= 16'h03cf;
        coeff[380] <= 16'h03d2;
        coeff[381] <= 16'h03d6;
        coeff[382] <= 16'h03d6;
        coeff[383] <= 16'h03d9;
        coeff[384] <= 16'h03dc;
        coeff[385] <= 16'h03dc;
        coeff[386] <= 16'h03e0;
        coeff[387] <= 16'h03e0;
        coeff[388] <= 16'h03e3;
        coeff[389] <= 16'h03e6;
        coeff[390] <= 16'h03e6;
        coeff[391] <= 16'h03e9;
        coeff[392] <= 16'h03ed;
        coeff[393] <= 16'h03ed;
        coeff[394] <= 16'h03f0;
        coeff[395] <= 16'h03f0;
        coeff[396] <= 16'h03f3;
        coeff[397] <= 16'h03f7;
        coeff[398] <= 16'h03f7;
        coeff[399] <= 16'h03fa;
        coeff[400] <= 16'h03fd;
        coeff[401] <= 16'h03fd;
        coeff[402] <= 16'h0400;
        coeff[403] <= 16'h0400;
        coeff[404] <= 16'h0404;
        coeff[405] <= 16'h0404;
        coeff[406] <= 16'h0407;
        coeff[407] <= 16'h040a;
        coeff[408] <= 16'h040a;
        coeff[409] <= 16'h040e;
        coeff[410] <= 16'h040e;
        coeff[411] <= 16'h0411;
        coeff[412] <= 16'h0414;
        coeff[413] <= 16'h0414;
        coeff[414] <= 16'h0418;
        coeff[415] <= 16'h0418;
        coeff[416] <= 16'h041b;
        coeff[417] <= 16'h041e;
        coeff[418] <= 16'h041e;
        coeff[419] <= 16'h0421;
        coeff[420] <= 16'h0421;
        coeff[421] <= 16'h0425;
        coeff[422] <= 16'h0428;
        coeff[423] <= 16'h0428;
        coeff[424] <= 16'h042b;
        coeff[425] <= 16'h042b;
        coeff[426] <= 16'h042f;
        coeff[427] <= 16'h0432;
        coeff[428] <= 16'h0432;
        coeff[429] <= 16'h0435;
        coeff[430] <= 16'h0438;
        coeff[431] <= 16'h0438;
        coeff[432] <= 16'h043c;
        coeff[433] <= 16'h043c;
        coeff[434] <= 16'h043f;
        coeff[435] <= 16'h0442;
        coeff[436] <= 16'h0442;
        coeff[437] <= 16'h0446;
        coeff[438] <= 16'h0449;
        coeff[439] <= 16'h044c;
        coeff[440] <= 16'h044c;
        coeff[441] <= 16'h0450;
        coeff[442] <= 16'h0453;
        coeff[443] <= 16'h0453;
        coeff[444] <= 16'h0456;
        coeff[445] <= 16'h0459;
        coeff[446] <= 16'h045d;
        coeff[447] <= 16'h045d;
        coeff[448] <= 16'h0460;
        coeff[449] <= 16'h0463;
        coeff[450] <= 16'h0467;
        coeff[451] <= 16'h0467;
        coeff[452] <= 16'h046a;
        coeff[453] <= 16'h046d;
        coeff[454] <= 16'h0470;
        coeff[455] <= 16'h0474;
        coeff[456] <= 16'h0477;
        coeff[457] <= 16'h0477;
        coeff[458] <= 16'h047a;
        coeff[459] <= 16'h047e;
        coeff[460] <= 16'h0481;
        coeff[461] <= 16'h0484;
        coeff[462] <= 16'h0488;
        coeff[463] <= 16'h048b;
        coeff[464] <= 16'h048e;
        coeff[465] <= 16'h0491;
        coeff[466] <= 16'h0495;
        coeff[467] <= 16'h0498;
        coeff[468] <= 16'h049b;
        coeff[469] <= 16'h049f;
        coeff[470] <= 16'h04a2;
        coeff[471] <= 16'h04a5;
        coeff[472] <= 16'h04a8;
        coeff[473] <= 16'h04ac;
        coeff[474] <= 16'h04af;
        coeff[475] <= 16'h04b2;
        coeff[476] <= 16'h04b6;
        coeff[477] <= 16'h04b9;
        coeff[478] <= 16'h04c0;
        coeff[479] <= 16'h04c3;
        coeff[480] <= 16'h04c6;
        coeff[481] <= 16'h04c9;
        coeff[482] <= 16'h04cd;
        coeff[483] <= 16'h04d3;
        coeff[484] <= 16'h04d7;
        coeff[485] <= 16'h04da;
        coeff[486] <= 16'h04dd;
        coeff[487] <= 16'h04e4;
        coeff[488] <= 16'h04e7;
        coeff[489] <= 16'h04ee;
        coeff[490] <= 16'h04f1;
        coeff[491] <= 16'h04f4;
        coeff[492] <= 16'h04fb;
        coeff[493] <= 16'h04fe;
        coeff[494] <= 16'h0505;
        coeff[495] <= 16'h0508;
        coeff[496] <= 16'h050f;
        coeff[497] <= 16'h0512;
        coeff[498] <= 16'h0519;
        coeff[499] <= 16'h051c;
        coeff[500] <= 16'h0522;
        coeff[501] <= 16'h0526;
        coeff[502] <= 16'h052c;
        coeff[503] <= 16'h0533;
        coeff[504] <= 16'h0536;
        coeff[505] <= 16'h053d;
        coeff[506] <= 16'h0543;
        coeff[507] <= 16'h0547;
        coeff[508] <= 16'h054d;
        coeff[509] <= 16'h0554;
        coeff[510] <= 16'h055a;
        coeff[511] <= 16'h0561;
        coeff[512] <= 16'h0568;
        coeff[513] <= 16'h056b;
        coeff[514] <= 16'h0571;
        coeff[515] <= 16'h0578;
        coeff[516] <= 16'h057f;
        coeff[517] <= 16'h0585;
        coeff[518] <= 16'h058c;
        coeff[519] <= 16'h0592;
        coeff[520] <= 16'h0599;
        coeff[521] <= 16'h059c;
        coeff[522] <= 16'h05a3;
        coeff[523] <= 16'h05a9;
        coeff[524] <= 16'h05b0;
        coeff[525] <= 16'h05b7;
        coeff[526] <= 16'h05bd;
        coeff[527] <= 16'h05c4;
        coeff[528] <= 16'h05ca;
        coeff[529] <= 16'h05d1;
        coeff[530] <= 16'h05d8;
        coeff[531] <= 16'h05de;
        coeff[532] <= 16'h05e5;
        coeff[533] <= 16'h05eb;
        coeff[534] <= 16'h05f2;
        coeff[535] <= 16'h05f9;
        coeff[536] <= 16'h05ff;
        coeff[537] <= 16'h0606;
        coeff[538] <= 16'h060c;
        coeff[539] <= 16'h0613;
        coeff[540] <= 16'h0619;
        coeff[541] <= 16'h0620;
        coeff[542] <= 16'h0627;
        coeff[543] <= 16'h062d;
        coeff[544] <= 16'h0634;
        coeff[545] <= 16'h063a;
        coeff[546] <= 16'h0641;
        coeff[547] <= 16'h0648;
        coeff[548] <= 16'h064e;
        coeff[549] <= 16'h0655;
        coeff[550] <= 16'h065f;
        coeff[551] <= 16'h0665;
        coeff[552] <= 16'h066c;
        coeff[553] <= 16'h0672;
        coeff[554] <= 16'h0679;
        coeff[555] <= 16'h0680;
        coeff[556] <= 16'h0689;
        coeff[557] <= 16'h0690;
        coeff[558] <= 16'h0697;
        coeff[559] <= 16'h069d;
        coeff[560] <= 16'h06a7;
        coeff[561] <= 16'h06ae;
        coeff[562] <= 16'h06b4;
        coeff[563] <= 16'h06be;
        coeff[564] <= 16'h06c5;
        coeff[565] <= 16'h06cb;
        coeff[566] <= 16'h06d5;
        coeff[567] <= 16'h06dc;
        coeff[568] <= 16'h06e6;
        coeff[569] <= 16'h06ec;
        coeff[570] <= 16'h06f6;
        coeff[571] <= 16'h06fd;
        coeff[572] <= 16'h0707;
        coeff[573] <= 16'h070d;
        coeff[574] <= 16'h0717;
        coeff[575] <= 16'h071e;
        coeff[576] <= 16'h0728;
        coeff[577] <= 16'h072e;
        coeff[578] <= 16'h0738;
        coeff[579] <= 16'h0742;
        coeff[580] <= 16'h0749;
        coeff[581] <= 16'h0752;
        coeff[582] <= 16'h075c;
        coeff[583] <= 16'h0763;
        coeff[584] <= 16'h076d;
        coeff[585] <= 16'h0777;
        coeff[586] <= 16'h0781;
        coeff[587] <= 16'h078a;
        coeff[588] <= 16'h0794;
        coeff[589] <= 16'h079b;
        coeff[590] <= 16'h07a5;
        coeff[591] <= 16'h07af;
        coeff[592] <= 16'h07b9;
        coeff[593] <= 16'h07c2;
        coeff[594] <= 16'h07cc;
        coeff[595] <= 16'h07d6;
        coeff[596] <= 16'h07e0;
        coeff[597] <= 16'h07ea;
        coeff[598] <= 16'h07f7;
        coeff[599] <= 16'h0801;
        coeff[600] <= 16'h080b;
        coeff[601] <= 16'h0815;
        coeff[602] <= 16'h081f;
        coeff[603] <= 16'h082c;
        coeff[604] <= 16'h0836;
        coeff[605] <= 16'h0840;
        coeff[606] <= 16'h084d;
        coeff[607] <= 16'h0857;
        coeff[608] <= 16'h0864;
        coeff[609] <= 16'h086e;
        coeff[610] <= 16'h0878;
        coeff[611] <= 16'h0885;
        coeff[612] <= 16'h0892;
        coeff[613] <= 16'h089c;
        coeff[614] <= 16'h08a9;
        coeff[615] <= 16'h08b3;
        coeff[616] <= 16'h08c0;
        coeff[617] <= 16'h08cd;
        coeff[618] <= 16'h08da;
        coeff[619] <= 16'h08e4;
        coeff[620] <= 16'h08f1;
        coeff[621] <= 16'h08ff;
        coeff[622] <= 16'h090c;
        coeff[623] <= 16'h0919;
        coeff[624] <= 16'h0926;
        coeff[625] <= 16'h0933;
        coeff[626] <= 16'h0941;
        coeff[627] <= 16'h094e;
        coeff[628] <= 16'h095b;
        coeff[629] <= 16'h0968;
        coeff[630] <= 16'h0975;
        coeff[631] <= 16'h0986;
        coeff[632] <= 16'h0993;
        coeff[633] <= 16'h09a0;
        coeff[634] <= 16'h09b1;
        coeff[635] <= 16'h09be;
        coeff[636] <= 16'h09cb;
        coeff[637] <= 16'h09db;
        coeff[638] <= 16'h09e9;
        coeff[639] <= 16'h09f9;
        coeff[640] <= 16'h0a09;
        coeff[641] <= 16'h0a17;
        coeff[642] <= 16'h0a27;
        coeff[643] <= 16'h0a34;
        coeff[644] <= 16'h0a45;
        coeff[645] <= 16'h0a55;
        coeff[646] <= 16'h0a66;
        coeff[647] <= 16'h0a76;
        coeff[648] <= 16'h0a83;
        coeff[649] <= 16'h0a94;
        coeff[650] <= 16'h0aa4;
        coeff[651] <= 16'h0ab5;
        coeff[652] <= 16'h0ac5;
        coeff[653] <= 16'h0ad6;
        coeff[654] <= 16'h0ae6;
        coeff[655] <= 16'h0af7;
        coeff[656] <= 16'h0b07;
        coeff[657] <= 16'h0b18;
        coeff[658] <= 16'h0b2b;
        coeff[659] <= 16'h0b3c;
        coeff[660] <= 16'h0b4c;
        coeff[661] <= 16'h0b5d;
        coeff[662] <= 16'h0b71;
        coeff[663] <= 16'h0b81;
        coeff[664] <= 16'h0b91;
        coeff[665] <= 16'h0ba5;
        coeff[666] <= 16'h0bb6;
        coeff[667] <= 16'h0bc6;
        coeff[668] <= 16'h0bda;
        coeff[669] <= 16'h0bea;
        coeff[670] <= 16'h0bfe;
        coeff[671] <= 16'h0c12;
        coeff[672] <= 16'h0c22;
        coeff[673] <= 16'h0c36;
        coeff[674] <= 16'h0c47;
        coeff[675] <= 16'h0c5a;
        coeff[676] <= 16'h0c6e;
        coeff[677] <= 16'h0c7f;
        coeff[678] <= 16'h0c92;
        coeff[679] <= 16'h0ca6;
        coeff[680] <= 16'h0cba;
        coeff[681] <= 16'h0cce;
        coeff[682] <= 16'h0ce1;
        coeff[683] <= 16'h0cf2;
        coeff[684] <= 16'h0d06;
        coeff[685] <= 16'h0d19;
        coeff[686] <= 16'h0d2d;
        coeff[687] <= 16'h0d41;
        coeff[688] <= 16'h0d55;
        coeff[689] <= 16'h0d69;
        coeff[690] <= 16'h0d7c;
        coeff[691] <= 16'h0d93;
        coeff[692] <= 16'h0da7;
        coeff[693] <= 16'h0dbb;
        coeff[694] <= 16'h0dcf;
        coeff[695] <= 16'h0de2;
        coeff[696] <= 16'h0df9;
        coeff[697] <= 16'h0e0d;
        coeff[698] <= 16'h0e21;
        coeff[699] <= 16'h0e38;
        coeff[700] <= 16'h0e4c;
        coeff[701] <= 16'h0e60;
        coeff[702] <= 16'h0e77;
        coeff[703] <= 16'h0e8a;
        coeff[704] <= 16'h0ea2;
        coeff[705] <= 16'h0eb5;
        coeff[706] <= 16'h0ecc;
        coeff[707] <= 16'h0ee0;
        coeff[708] <= 16'h0ef7;
        coeff[709] <= 16'h0f0b;
        coeff[710] <= 16'h0f22;
        coeff[711] <= 16'h0f39;
        coeff[712] <= 16'h0f4d;
        coeff[713] <= 16'h0f64;
        coeff[714] <= 16'h0f7b;
        coeff[715] <= 16'h0f8f;
        coeff[716] <= 16'h0fa6;
        coeff[717] <= 16'h0fbd;
        coeff[718] <= 16'h0fd4;
        coeff[719] <= 16'h0feb;
        coeff[720] <= 16'h0fff;
        coeff[721] <= 16'h1016;
        coeff[722] <= 16'h102d;
        coeff[723] <= 16'h1044;
        coeff[724] <= 16'h105b;
        coeff[725] <= 16'h1072;
        coeff[726] <= 16'h1089;
        coeff[727] <= 16'h10a0;
        coeff[728] <= 16'h10b7;
        coeff[729] <= 16'h10ce;
        coeff[730] <= 16'h10e5;
        coeff[731] <= 16'h1100;
        coeff[732] <= 16'h1117;
        coeff[733] <= 16'h112e;
        coeff[734] <= 16'h1145;
        coeff[735] <= 16'h115c;
        coeff[736] <= 16'h1176;
        coeff[737] <= 16'h118d;
        coeff[738] <= 16'h11a4;
        coeff[739] <= 16'h11bb;
        coeff[740] <= 16'h11d6;
        coeff[741] <= 16'h11ed;
        coeff[742] <= 16'h1204;
        coeff[743] <= 16'h121e;
        coeff[744] <= 16'h1235;
        coeff[745] <= 16'h1250;
        coeff[746] <= 16'h1267;
        coeff[747] <= 16'h1281;
        coeff[748] <= 16'h1298;
        coeff[749] <= 16'h12b2;
        coeff[750] <= 16'h12ca;
        coeff[751] <= 16'h12e4;
        coeff[752] <= 16'h12fb;
        coeff[753] <= 16'h1315;
        coeff[754] <= 16'h1330;
        coeff[755] <= 16'h1347;
        coeff[756] <= 16'h1361;
        coeff[757] <= 16'h137b;
        coeff[758] <= 16'h1392;
        coeff[759] <= 16'h13ad;
        coeff[760] <= 16'h13c7;
        coeff[761] <= 16'h13e2;
        coeff[762] <= 16'h13f9;
        coeff[763] <= 16'h1413;
        coeff[764] <= 16'h142d;
        coeff[765] <= 16'h1448;
        coeff[766] <= 16'h1462;
        coeff[767] <= 16'h147c;
        coeff[768] <= 16'h1497;
        coeff[769] <= 16'h14ae;
        coeff[770] <= 16'h14cb;
        coeff[771] <= 16'h14e6;
        coeff[772] <= 16'h1500;
        coeff[773] <= 16'h151e;
        coeff[774] <= 16'h1538;
        coeff[775] <= 16'h1556;
        coeff[776] <= 16'h1573;
        coeff[777] <= 16'h1591;
        coeff[778] <= 16'h15af;
        coeff[779] <= 16'h15d0;
        coeff[780] <= 16'h15ed;
        coeff[781] <= 16'h160b;
        coeff[782] <= 16'h162c;
        coeff[783] <= 16'h164d;
        coeff[784] <= 16'h166e;
        coeff[785] <= 16'h168f;
        coeff[786] <= 16'h16b0;
        coeff[787] <= 16'h16d1;
        coeff[788] <= 16'h16f2;
        coeff[789] <= 16'h1712;
        coeff[790] <= 16'h1737;
        coeff[791] <= 16'h1758;
        coeff[792] <= 16'h177c;
        coeff[793] <= 16'h17a0;
        coeff[794] <= 16'h17c1;
        coeff[795] <= 16'h17e5;
        coeff[796] <= 16'h180a;
        coeff[797] <= 16'h182e;
        coeff[798] <= 16'h1852;
        coeff[799] <= 16'h187a;
        coeff[800] <= 16'h189e;
        coeff[801] <= 16'h18c2;
        coeff[802] <= 16'h18ea;
        coeff[803] <= 16'h190e;
        coeff[804] <= 16'h1935;
        coeff[805] <= 16'h195a;
        coeff[806] <= 16'h1981;
        coeff[807] <= 16'h19a9;
        coeff[808] <= 16'h19cd;
        coeff[809] <= 16'h19f4;
        coeff[810] <= 16'h1a1c;
        coeff[811] <= 16'h1a43;
        coeff[812] <= 16'h1a6b;
        coeff[813] <= 16'h1a93;
        coeff[814] <= 16'h1aba;
        coeff[815] <= 16'h1ae2;
        coeff[816] <= 16'h1b09;
        coeff[817] <= 16'h1b34;
        coeff[818] <= 16'h1b5b;
        coeff[819] <= 16'h1b83;
        coeff[820] <= 16'h1bab;
        coeff[821] <= 16'h1bd5;
        coeff[822] <= 16'h1bfd;
        coeff[823] <= 16'h1c24;
        coeff[824] <= 16'h1c4f;
        coeff[825] <= 16'h1c77;
        coeff[826] <= 16'h1ca2;
        coeff[827] <= 16'h1cc9;
        coeff[828] <= 16'h1cf4;
        coeff[829] <= 16'h1d1b;
        coeff[830] <= 16'h1d46;
        coeff[831] <= 16'h1d6e;
        coeff[832] <= 16'h1d99;
        coeff[833] <= 16'h1dc0;
        coeff[834] <= 16'h1deb;
        coeff[835] <= 16'h1e13;
        coeff[836] <= 16'h1e3d;
        coeff[837] <= 16'h1e68;
        coeff[838] <= 16'h1e90;
        coeff[839] <= 16'h1ebb;
        coeff[840] <= 16'h1ee5;
        coeff[841] <= 16'h1f10;
        coeff[842] <= 16'h1f3b;
        coeff[843] <= 16'h1f66;
        coeff[844] <= 16'h1f91;
        coeff[845] <= 16'h1fbb;
        coeff[846] <= 16'h1fe6;
        coeff[847] <= 16'h2011;
        coeff[848] <= 16'h203f;
        coeff[849] <= 16'h206a;
        coeff[850] <= 16'h2095;
        coeff[851] <= 16'h20c3;
        coeff[852] <= 16'h20ee;
        coeff[853] <= 16'h211c;
        coeff[854] <= 16'h2147;
        coeff[855] <= 16'h2175;
        coeff[856] <= 16'h21a3;
        coeff[857] <= 16'h21ce;
        coeff[858] <= 16'h21fc;
        coeff[859] <= 16'h222a;
        coeff[860] <= 16'h2258;
        coeff[861] <= 16'h2286;
        coeff[862] <= 16'h22b1;
        coeff[863] <= 16'h22df;
        coeff[864] <= 16'h2311;
        coeff[865] <= 16'h233f;
        coeff[866] <= 16'h236d;
        coeff[867] <= 16'h239b;
        coeff[868] <= 16'h23c9;
        coeff[869] <= 16'h23f7;
        coeff[870] <= 16'h2429;
        coeff[871] <= 16'h2457;
        coeff[872] <= 16'h2488;
        coeff[873] <= 16'h24b6;
        coeff[874] <= 16'h24e8;
        coeff[875] <= 16'h2516;
        coeff[876] <= 16'h2547;
        coeff[877] <= 16'h2575;
        coeff[878] <= 16'h25a7;
        coeff[879] <= 16'h25d8;
        coeff[880] <= 16'h260a;
        coeff[881] <= 16'h263b;
        coeff[882] <= 16'h266c;
        coeff[883] <= 16'h269e;
        coeff[884] <= 16'h26cf;
        coeff[885] <= 16'h2701;
        coeff[886] <= 16'h2732;
        coeff[887] <= 16'h2764;
        coeff[888] <= 16'h2795;
        coeff[889] <= 16'h27c6;
        coeff[890] <= 16'h27fb;
        coeff[891] <= 16'h282c;
        coeff[892] <= 16'h285e;
        coeff[893] <= 16'h2893;
        coeff[894] <= 16'h28c4;
        coeff[895] <= 16'h28f9;
        coeff[896] <= 16'h292d;
        coeff[897] <= 16'h295f;
        coeff[898] <= 16'h2994;
        coeff[899] <= 16'h29c8;
        coeff[900] <= 16'h29fa;
        coeff[901] <= 16'h2a2e;
        coeff[902] <= 16'h2a63;
        coeff[903] <= 16'h2a98;
        coeff[904] <= 16'h2acd;
        coeff[905] <= 16'h2b01;
        coeff[906] <= 16'h2b36;
        coeff[907] <= 16'h2b6b;
        coeff[908] <= 16'h2ba3;
        coeff[909] <= 16'h2bd7;
        coeff[910] <= 16'h2c0c;
        coeff[911] <= 16'h2c41;
        coeff[912] <= 16'h2c79;
        coeff[913] <= 16'h2cad;
        coeff[914] <= 16'h2ce5;
        coeff[915] <= 16'h2d1a;
        coeff[916] <= 16'h2d52;
        coeff[917] <= 16'h2d87;
        coeff[918] <= 16'h2dbf;
        coeff[919] <= 16'h2df7;
        coeff[920] <= 16'h2e2f;
        coeff[921] <= 16'h2e64;
        coeff[922] <= 16'h2e9c;
        coeff[923] <= 16'h2ed4;
        coeff[924] <= 16'h2f0c;
        coeff[925] <= 16'h2f44;
        coeff[926] <= 16'h2f7c;
        coeff[927] <= 16'h2fb4;
        coeff[928] <= 16'h2fef;
        coeff[929] <= 16'h3027;
        coeff[930] <= 16'h305f;
        coeff[931] <= 16'h3097;
        coeff[932] <= 16'h30d2;
        coeff[933] <= 16'h310a;
        coeff[934] <= 16'h3145;
        coeff[935] <= 16'h317d;
        coeff[936] <= 16'h31b9;
        coeff[937] <= 16'h31f1;
        coeff[938] <= 16'h322c;
        coeff[939] <= 16'h3267;
        coeff[940] <= 16'h329f;
        coeff[941] <= 16'h32db;
        coeff[942] <= 16'h3316;
        coeff[943] <= 16'h3351;
        coeff[944] <= 16'h338d;
        coeff[945] <= 16'h33c8;
        coeff[946] <= 16'h3403;
        coeff[947] <= 16'h343e;
        coeff[948] <= 16'h347a;
        coeff[949] <= 16'h34b5;
        coeff[950] <= 16'h34f0;
        coeff[951] <= 16'h352f;
        coeff[952] <= 16'h356a;
        coeff[953] <= 16'h35a6;
        coeff[954] <= 16'h35e4;
        coeff[955] <= 16'h361f;
        coeff[956] <= 16'h365e;
        coeff[957] <= 16'h3699;
        coeff[958] <= 16'h36d8;
        coeff[959] <= 16'h3716;
        coeff[960] <= 16'h3755;
        coeff[961] <= 16'h3790;
        coeff[962] <= 16'h37d2;
        coeff[963] <= 16'h3811;
        coeff[964] <= 16'h3853;
        coeff[965] <= 16'h3895;
        coeff[966] <= 16'h38d6;
        coeff[967] <= 16'h391c;
        coeff[968] <= 16'h3961;
        coeff[969] <= 16'h39a6;
        coeff[970] <= 16'h39eb;
        coeff[971] <= 16'h3a34;
        coeff[972] <= 16'h3a79;
        coeff[973] <= 16'h3ac1;
        coeff[974] <= 16'h3b0a;
        coeff[975] <= 16'h3b56;
        coeff[976] <= 16'h3b9e;
        coeff[977] <= 16'h3be6;
        coeff[978] <= 16'h3c32;
        coeff[979] <= 16'h3c7e;
        coeff[980] <= 16'h3cc7;
        coeff[981] <= 16'h3d12;
        coeff[982] <= 16'h3d5e;
        coeff[983] <= 16'h3daa;
        coeff[984] <= 16'h3df6;
        coeff[985] <= 16'h3e41;
        coeff[986] <= 16'h3e8d;
        coeff[987] <= 16'h3ed9;
        coeff[988] <= 16'h3f25;
        coeff[989] <= 16'h3f74;
        coeff[990] <= 16'h3fbf;
        coeff[991] <= 16'h400b;
        coeff[992] <= 16'h4057;
        coeff[993] <= 16'h409f;
        coeff[994] <= 16'h40eb;
        coeff[995] <= 16'h4137;
        coeff[996] <= 16'h4186;
        coeff[997] <= 16'h41d2;
        coeff[998] <= 16'h4221;
        coeff[999] <= 16'h4270;
        coeff[1000] <= 16'h42bf;
        coeff[1001] <= 16'h4311;
        coeff[1002] <= 16'h4364;
        coeff[1003] <= 16'h43b6;
        coeff[1004] <= 16'h440f;
        coeff[1005] <= 16'h4465;
        coeff[1006] <= 16'h44c1;
        coeff[1007] <= 16'h451d;
        coeff[1008] <= 16'h457d;
        coeff[1009] <= 16'h45df;
        coeff[1010] <= 16'h4650;
        coeff[1011] <= 16'h46c6;
        coeff[1012] <= 16'h4747;
        coeff[1013] <= 16'h47c7;
        coeff[1014] <= 16'h484e;
        coeff[1015] <= 16'h48d2;
        coeff[1016] <= 16'h4959;
        coeff[1017] <= 16'h49dd;
        coeff[1018] <= 16'h4a67;
        coeff[1019] <= 16'h4af1;
        coeff[1020] <= 16'h4b7f;
        coeff[1021] <= 16'h4c10;
        coeff[1022] <= 16'h4ca1;
        coeff[1023] <= 16'h4d35;
        coeff[1024] <= 16'h3b31;
        coeff[1025] <= 16'h3b87;
        coeff[1026] <= 16'h3bdd;
        coeff[1027] <= 16'h3c36;
        coeff[1028] <= 16'h3c88;
        coeff[1029] <= 16'h3cda;
        coeff[1030] <= 16'h3d2d;
        coeff[1031] <= 16'h3d78;
        coeff[1032] <= 16'h3dc4;
        coeff[1033] <= 16'h3e09;
        coeff[1034] <= 16'h3e52;
        coeff[1035] <= 16'h3e97;
        coeff[1036] <= 16'h3edc;
        coeff[1037] <= 16'h3f21;
        coeff[1038] <= 16'h3f67;
        coeff[1039] <= 16'h3fac;
        coeff[1040] <= 16'h3ff1;
        coeff[1041] <= 16'h4033;
        coeff[1042] <= 16'h4078;
        coeff[1043] <= 16'h40ba;
        coeff[1044] <= 16'h40ff;
        coeff[1045] <= 16'h4141;
        coeff[1046] <= 16'h4186;
        coeff[1047] <= 16'h41c8;
        coeff[1048] <= 16'h420d;
        coeff[1049] <= 16'h424f;
        coeff[1050] <= 16'h4294;
        coeff[1051] <= 16'h42d6;
        coeff[1052] <= 16'h431b;
        coeff[1053] <= 16'h4360;
        coeff[1054] <= 16'h43a6;
        coeff[1055] <= 16'h43eb;
        coeff[1056] <= 16'h4433;
        coeff[1057] <= 16'h4478;
        coeff[1058] <= 16'h44c1;
        coeff[1059] <= 16'h4506;
        coeff[1060] <= 16'h454f;
        coeff[1061] <= 16'h4597;
        coeff[1062] <= 16'h45df;
        coeff[1063] <= 16'h462b;
        coeff[1064] <= 16'h4674;
        coeff[1065] <= 16'h46bc;
        coeff[1066] <= 16'h4705;
        coeff[1067] <= 16'h4750;
        coeff[1068] <= 16'h4799;
        coeff[1069] <= 16'h47e5;
        coeff[1070] <= 16'h482d;
        coeff[1071] <= 16'h4879;
        coeff[1072] <= 16'h48c1;
        coeff[1073] <= 16'h490a;
        coeff[1074] <= 16'h4956;
        coeff[1075] <= 16'h499e;
        coeff[1076] <= 16'h49e7;
        coeff[1077] <= 16'h4a2f;
        coeff[1078] <= 16'h4a78;
        coeff[1079] <= 16'h4ac0;
        coeff[1080] <= 16'h4b08;
        coeff[1081] <= 16'h4b51;
        coeff[1082] <= 16'h4b96;
        coeff[1083] <= 16'h4bdb;
        coeff[1084] <= 16'h4c24;
        coeff[1085] <= 16'h4c69;
        coeff[1086] <= 16'h4cab;
        coeff[1087] <= 16'h4cf0;
        coeff[1088] <= 16'h4d35;
        coeff[1089] <= 16'h4d77;
        coeff[1090] <= 16'h4db9;
        coeff[1091] <= 16'h4dfb;
        coeff[1092] <= 16'h4e39;
        coeff[1093] <= 16'h4e7b;
        coeff[1094] <= 16'h4eba;
        coeff[1095] <= 16'h4ef8;
        coeff[1096] <= 16'h4f3a;
        coeff[1097] <= 16'h4f79;
        coeff[1098] <= 16'h4fb4;
        coeff[1099] <= 16'h4ff3;
        coeff[1100] <= 16'h5031;
        coeff[1101] <= 16'h506d;
        coeff[1102] <= 16'h50ab;
        coeff[1103] <= 16'h50e7;
        coeff[1104] <= 16'h5125;
        coeff[1105] <= 16'h5161;
        coeff[1106] <= 16'h519c;
        coeff[1107] <= 16'h51da;
        coeff[1108] <= 16'h5216;
        coeff[1109] <= 16'h5251;
        coeff[1110] <= 16'h528c;
        coeff[1111] <= 16'h52cb;
        coeff[1112] <= 16'h5306;
        coeff[1113] <= 16'h5341;
        coeff[1114] <= 16'h537d;
        coeff[1115] <= 16'h53bb;
        coeff[1116] <= 16'h53f7;
        coeff[1117] <= 16'h5435;
        coeff[1118] <= 16'h5471;
        coeff[1119] <= 16'h54af;
        coeff[1120] <= 16'h54ee;
        coeff[1121] <= 16'h5529;
        coeff[1122] <= 16'h5568;
        coeff[1123] <= 16'h55a6;
        coeff[1124] <= 16'h55e5;
        coeff[1125] <= 16'h5623;
        coeff[1126] <= 16'h5662;
        coeff[1127] <= 16'h569d;
        coeff[1128] <= 16'h56dc;
        coeff[1129] <= 16'h571a;
        coeff[1130] <= 16'h5759;
        coeff[1131] <= 16'h5798;
        coeff[1132] <= 16'h57d6;
        coeff[1133] <= 16'h5815;
        coeff[1134] <= 16'h5853;
        coeff[1135] <= 16'h5892;
        coeff[1136] <= 16'h58d1;
        coeff[1137] <= 16'h590f;
        coeff[1138] <= 16'h594e;
        coeff[1139] <= 16'h598c;
        coeff[1140] <= 16'h59c8;
        coeff[1141] <= 16'h5a06;
        coeff[1142] <= 16'h5a45;
        coeff[1143] <= 16'h5a83;
        coeff[1144] <= 16'h5abf;
        coeff[1145] <= 16'h5afd;
        coeff[1146] <= 16'h5b39;
        coeff[1147] <= 16'h5b77;
        coeff[1148] <= 16'h5bb2;
        coeff[1149] <= 16'h5bf1;
        coeff[1150] <= 16'h5c2c;
        coeff[1151] <= 16'h5c68;
        coeff[1152] <= 16'h5ca6;
        coeff[1153] <= 16'h5ce2;
        coeff[1154] <= 16'h5d1d;
        coeff[1155] <= 16'h5d58;
        coeff[1156] <= 16'h5d93;
        coeff[1157] <= 16'h5dcf;
        coeff[1158] <= 16'h5e0a;
        coeff[1159] <= 16'h5e45;
        coeff[1160] <= 16'h5e81;
        coeff[1161] <= 16'h5ebc;
        coeff[1162] <= 16'h5ef7;
        coeff[1163] <= 16'h5f32;
        coeff[1164] <= 16'h5f6e;
        coeff[1165] <= 16'h5fa9;
        coeff[1166] <= 16'h5fe4;
        coeff[1167] <= 16'h6020;
        coeff[1168] <= 16'h605b;
        coeff[1169] <= 16'h6093;
        coeff[1170] <= 16'h60ce;
        coeff[1171] <= 16'h610a;
        coeff[1172] <= 16'h6145;
        coeff[1173] <= 16'h6180;
        coeff[1174] <= 16'h61bb;
        coeff[1175] <= 16'h61f7;
        coeff[1176] <= 16'h622f;
        coeff[1177] <= 16'h626a;
        coeff[1178] <= 16'h62a5;
        coeff[1179] <= 16'h62e1;
        coeff[1180] <= 16'h631c;
        coeff[1181] <= 16'h6354;
        coeff[1182] <= 16'h638f;
        coeff[1183] <= 16'h63cb;
        coeff[1184] <= 16'h6406;
        coeff[1185] <= 16'h643e;
        coeff[1186] <= 16'h6479;
        coeff[1187] <= 16'h64b4;
        coeff[1188] <= 16'h64f0;
        coeff[1189] <= 16'h6528;
        coeff[1190] <= 16'h6563;
        coeff[1191] <= 16'h659e;
        coeff[1192] <= 16'h65d6;
        coeff[1193] <= 16'h6612;
        coeff[1194] <= 16'h664d;
        coeff[1195] <= 16'h6688;
        coeff[1196] <= 16'h66c0;
        coeff[1197] <= 16'h66fb;
        coeff[1198] <= 16'h6737;
        coeff[1199] <= 16'h676f;
        coeff[1200] <= 16'h67aa;
        coeff[1201] <= 16'h67e5;
        coeff[1202] <= 16'h6821;
        coeff[1203] <= 16'h6859;
        coeff[1204] <= 16'h6894;
        coeff[1205] <= 16'h68cf;
        coeff[1206] <= 16'h6907;
        coeff[1207] <= 16'h6943;
        coeff[1208] <= 16'h697e;
        coeff[1209] <= 16'h69b6;
        coeff[1210] <= 16'h69f1;
        coeff[1211] <= 16'h6a2c;
        coeff[1212] <= 16'h6a68;
        coeff[1213] <= 16'h6aa0;
        coeff[1214] <= 16'h6adb;
        coeff[1215] <= 16'h6b16;
        coeff[1216] <= 16'h6b52;
        coeff[1217] <= 16'h6b8a;
        coeff[1218] <= 16'h6bc5;
        coeff[1219] <= 16'h6c00;
        coeff[1220] <= 16'h6c38;
        coeff[1221] <= 16'h6c74;
        coeff[1222] <= 16'h6caf;
        coeff[1223] <= 16'h6cea;
        coeff[1224] <= 16'h6d25;
        coeff[1225] <= 16'h6d5d;
        coeff[1226] <= 16'h6d99;
        coeff[1227] <= 16'h6dd4;
        coeff[1228] <= 16'h6e0f;
        coeff[1229] <= 16'h6e4b;
        coeff[1230] <= 16'h6e83;
        coeff[1231] <= 16'h6ebe;
        coeff[1232] <= 16'h6ef9;
        coeff[1233] <= 16'h6f34;
        coeff[1234] <= 16'h6f70;
        coeff[1235] <= 16'h6fab;
        coeff[1236] <= 16'h6fe6;
        coeff[1237] <= 16'h7022;
        coeff[1238] <= 16'h705a;
        coeff[1239] <= 16'h7095;
        coeff[1240] <= 16'h70d0;
        coeff[1241] <= 16'h710c;
        coeff[1242] <= 16'h7147;
        coeff[1243] <= 16'h7182;
        coeff[1244] <= 16'h71bd;
        coeff[1245] <= 16'h71f9;
        coeff[1246] <= 16'h7234;
        coeff[1247] <= 16'h726f;
        coeff[1248] <= 16'h72ab;
        coeff[1249] <= 16'h72e6;
        coeff[1250] <= 16'h7324;
        coeff[1251] <= 16'h7360;
        coeff[1252] <= 16'h739b;
        coeff[1253] <= 16'h73d6;
        coeff[1254] <= 16'h7412;
        coeff[1255] <= 16'h744d;
        coeff[1256] <= 16'h7488;
        coeff[1257] <= 16'h74c7;
        coeff[1258] <= 16'h7502;
        coeff[1259] <= 16'h753d;
        coeff[1260] <= 16'h7579;
        coeff[1261] <= 16'h75b7;
        coeff[1262] <= 16'h75f3;
        coeff[1263] <= 16'h762e;
        coeff[1264] <= 16'h766d;
        coeff[1265] <= 16'h76a8;
        coeff[1266] <= 16'h76e3;
        coeff[1267] <= 16'h7722;
        coeff[1268] <= 16'h775d;
        coeff[1269] <= 16'h779c;
        coeff[1270] <= 16'h77d7;
        coeff[1271] <= 16'h7815;
        coeff[1272] <= 16'h7851;
        coeff[1273] <= 16'h788f;
        coeff[1274] <= 16'h78cb;
        coeff[1275] <= 16'h7909;
        coeff[1276] <= 16'h7948;
        coeff[1277] <= 16'h7983;
        coeff[1278] <= 16'h79c2;
        coeff[1279] <= 16'h7a00;
        coeff[1280] <= 16'h7a3f;
        coeff[1281] <= 16'h7a7a;
        coeff[1282] <= 16'h7ab9;
        coeff[1283] <= 16'h7af7;
        coeff[1284] <= 16'h7b36;
        coeff[1285] <= 16'h7b75;
        coeff[1286] <= 16'h7bb0;
        coeff[1287] <= 16'h7bee;
        coeff[1288] <= 16'h7c2d;
        coeff[1289] <= 16'h7c6c;
        coeff[1290] <= 16'h7caa;
        coeff[1291] <= 16'h7ce9;
        coeff[1292] <= 16'h7d27;
        coeff[1293] <= 16'h7d66;
        coeff[1294] <= 16'h7da5;
        coeff[1295] <= 16'h7de3;
        coeff[1296] <= 16'h7e22;
        coeff[1297] <= 16'h7e64;
        coeff[1298] <= 16'h7ea2;
        coeff[1299] <= 16'h7ee1;
        coeff[1300] <= 16'h7f1f;
        coeff[1301] <= 16'h7f5e;
        coeff[1302] <= 16'h7f9d;
        coeff[1303] <= 16'h7fde;
        coeff[1304] <= 16'h801d;
        coeff[1305] <= 16'h805c;
        coeff[1306] <= 16'h809a;
        coeff[1307] <= 16'h80dc;
        coeff[1308] <= 16'h811b;
        coeff[1309] <= 16'h8159;
        coeff[1310] <= 16'h819b;
        coeff[1311] <= 16'h81da;
        coeff[1312] <= 16'h8218;
        coeff[1313] <= 16'h825a;
        coeff[1314] <= 16'h8299;
        coeff[1315] <= 16'h82db;
        coeff[1316] <= 16'h8319;
        coeff[1317] <= 16'h835b;
        coeff[1318] <= 16'h839a;
        coeff[1319] <= 16'h83d8;
        coeff[1320] <= 16'h841a;
        coeff[1321] <= 16'h8459;
        coeff[1322] <= 16'h849b;
        coeff[1323] <= 16'h84dd;
        coeff[1324] <= 16'h851b;
        coeff[1325] <= 16'h855d;
        coeff[1326] <= 16'h859c;
        coeff[1327] <= 16'h85de;
        coeff[1328] <= 16'h861c;
        coeff[1329] <= 16'h865e;
        coeff[1330] <= 16'h86a0;
        coeff[1331] <= 16'h86de;
        coeff[1332] <= 16'h8720;
        coeff[1333] <= 16'h875f;
        coeff[1334] <= 16'h87a1;
        coeff[1335] <= 16'h87e3;
        coeff[1336] <= 16'h8821;
        coeff[1337] <= 16'h8863;
        coeff[1338] <= 16'h88a5;
        coeff[1339] <= 16'h88e4;
        coeff[1340] <= 16'h8926;
        coeff[1341] <= 16'h8967;
        coeff[1342] <= 16'h89a9;
        coeff[1343] <= 16'h89e8;
        coeff[1344] <= 16'h8a2a;
        coeff[1345] <= 16'h8a6c;
        coeff[1346] <= 16'h8aaa;
        coeff[1347] <= 16'h8aec;
        coeff[1348] <= 16'h8b2e;
        coeff[1349] <= 16'h8b70;
        coeff[1350] <= 16'h8baf;
        coeff[1351] <= 16'h8bf0;
        coeff[1352] <= 16'h8c32;
        coeff[1353] <= 16'h8c74;
        coeff[1354] <= 16'h8cb6;
        coeff[1355] <= 16'h8cf5;
        coeff[1356] <= 16'h8d37;
        coeff[1357] <= 16'h8d78;
        coeff[1358] <= 16'h8dba;
        coeff[1359] <= 16'h8df9;
        coeff[1360] <= 16'h8e3b;
        coeff[1361] <= 16'h8e7d;
        coeff[1362] <= 16'h8ebf;
        coeff[1363] <= 16'h8f00;
        coeff[1364] <= 16'h8f3f;
        coeff[1365] <= 16'h8f81;
        coeff[1366] <= 16'h8fc3;
        coeff[1367] <= 16'h9005;
        coeff[1368] <= 16'h9047;
        coeff[1369] <= 16'h9085;
        coeff[1370] <= 16'h90c7;
        coeff[1371] <= 16'h9109;
        coeff[1372] <= 16'h914b;
        coeff[1373] <= 16'h9189;
        coeff[1374] <= 16'h91cb;
        coeff[1375] <= 16'h920d;
        coeff[1376] <= 16'h924f;
        coeff[1377] <= 16'h9291;
        coeff[1378] <= 16'h92d0;
        coeff[1379] <= 16'h9311;
        coeff[1380] <= 16'h9353;
        coeff[1381] <= 16'h9395;
        coeff[1382] <= 16'h93d4;
        coeff[1383] <= 16'h9416;
        coeff[1384] <= 16'h9458;
        coeff[1385] <= 16'h9499;
        coeff[1386] <= 16'h94d8;
        coeff[1387] <= 16'h951a;
        coeff[1388] <= 16'h955c;
        coeff[1389] <= 16'h959e;
        coeff[1390] <= 16'h95dc;
        coeff[1391] <= 16'h961e;
        coeff[1392] <= 16'h9660;
        coeff[1393] <= 16'h969f;
        coeff[1394] <= 16'h96e0;
        coeff[1395] <= 16'h9722;
        coeff[1396] <= 16'h9761;
        coeff[1397] <= 16'h97a3;
        coeff[1398] <= 16'h97e5;
        coeff[1399] <= 16'h9823;
        coeff[1400] <= 16'h9865;
        coeff[1401] <= 16'h98a4;
        coeff[1402] <= 16'h98e6;
        coeff[1403] <= 16'h9928;
        coeff[1404] <= 16'h9966;
        coeff[1405] <= 16'h99a8;
        coeff[1406] <= 16'h99e7;
        coeff[1407] <= 16'h9a28;
        coeff[1408] <= 16'h9a6a;
        coeff[1409] <= 16'h9aa9;
        coeff[1410] <= 16'h9aeb;
        coeff[1411] <= 16'h9b29;
        coeff[1412] <= 16'h9b6b;
        coeff[1413] <= 16'h9bad;
        coeff[1414] <= 16'h9bef;
        coeff[1415] <= 16'h9c31;
        coeff[1416] <= 16'h9c73;
        coeff[1417] <= 16'h9cb5;
        coeff[1418] <= 16'h9cf7;
        coeff[1419] <= 16'h9d39;
        coeff[1420] <= 16'h9d7a;
        coeff[1421] <= 16'h9dbc;
        coeff[1422] <= 16'h9dfe;
        coeff[1423] <= 16'h9e43;
        coeff[1424] <= 16'h9e85;
        coeff[1425] <= 16'h9ec7;
        coeff[1426] <= 16'h9f0c;
        coeff[1427] <= 16'h9f4e;
        coeff[1428] <= 16'h9f90;
        coeff[1429] <= 16'h9fd5;
        coeff[1430] <= 16'ha017;
        coeff[1431] <= 16'ha05c;
        coeff[1432] <= 16'ha0a1;
        coeff[1433] <= 16'ha0e3;
        coeff[1434] <= 16'ha129;
        coeff[1435] <= 16'ha16a;
        coeff[1436] <= 16'ha1b0;
        coeff[1437] <= 16'ha1f5;
        coeff[1438] <= 16'ha237;
        coeff[1439] <= 16'ha27c;
        coeff[1440] <= 16'ha2c1;
        coeff[1441] <= 16'ha306;
        coeff[1442] <= 16'ha348;
        coeff[1443] <= 16'ha38d;
        coeff[1444] <= 16'ha3d2;
        coeff[1445] <= 16'ha418;
        coeff[1446] <= 16'ha45d;
        coeff[1447] <= 16'ha49f;
        coeff[1448] <= 16'ha4e4;
        coeff[1449] <= 16'ha529;
        coeff[1450] <= 16'ha56e;
        coeff[1451] <= 16'ha5b3;
        coeff[1452] <= 16'ha5f9;
        coeff[1453] <= 16'ha63a;
        coeff[1454] <= 16'ha680;
        coeff[1455] <= 16'ha6c5;
        coeff[1456] <= 16'ha70a;
        coeff[1457] <= 16'ha74f;
        coeff[1458] <= 16'ha794;
        coeff[1459] <= 16'ha7d6;
        coeff[1460] <= 16'ha81b;
        coeff[1461] <= 16'ha861;
        coeff[1462] <= 16'ha8a6;
        coeff[1463] <= 16'ha8e8;
        coeff[1464] <= 16'ha92d;
        coeff[1465] <= 16'ha972;
        coeff[1466] <= 16'ha9b4;
        coeff[1467] <= 16'ha9f9;
        coeff[1468] <= 16'haa3e;
        coeff[1469] <= 16'haa80;
        coeff[1470] <= 16'haac5;
        coeff[1471] <= 16'hab07;
        coeff[1472] <= 16'hab4c;
        coeff[1473] <= 16'hab8e;
        coeff[1474] <= 16'habd3;
        coeff[1475] <= 16'hac15;
        coeff[1476] <= 16'hac5a;
        coeff[1477] <= 16'hac9c;
        coeff[1478] <= 16'hacde;
        coeff[1479] <= 16'had23;
        coeff[1480] <= 16'had65;
        coeff[1481] <= 16'hada7;
        coeff[1482] <= 16'hade9;
        coeff[1483] <= 16'hae2b;
        coeff[1484] <= 16'hae6d;
        coeff[1485] <= 16'haeaf;
        coeff[1486] <= 16'haef1;
        coeff[1487] <= 16'haf33;
        coeff[1488] <= 16'haf74;
        coeff[1489] <= 16'hafb6;
        coeff[1490] <= 16'haff8;
        coeff[1491] <= 16'hb03a;
        coeff[1492] <= 16'hb079;
        coeff[1493] <= 16'hb0bb;
        coeff[1494] <= 16'hb0f9;
        coeff[1495] <= 16'hb13b;
        coeff[1496] <= 16'hb17a;
        coeff[1497] <= 16'hb1b8;
        coeff[1498] <= 16'hb1fa;
        coeff[1499] <= 16'hb239;
        coeff[1500] <= 16'hb277;
        coeff[1501] <= 16'hb2b6;
        coeff[1502] <= 16'hb2f4;
        coeff[1503] <= 16'hb333;
        coeff[1504] <= 16'hb372;
        coeff[1505] <= 16'hb3b0;
        coeff[1506] <= 16'hb3eb;
        coeff[1507] <= 16'hb42a;
        coeff[1508] <= 16'hb465;
        coeff[1509] <= 16'hb4a4;
        coeff[1510] <= 16'hb4df;
        coeff[1511] <= 16'hb51b;
        coeff[1512] <= 16'hb559;
        coeff[1513] <= 16'hb594;
        coeff[1514] <= 16'hb5d0;
        coeff[1515] <= 16'hb60b;
        coeff[1516] <= 16'hb643;
        coeff[1517] <= 16'hb67e;
        coeff[1518] <= 16'hb6ba;
        coeff[1519] <= 16'hb6f2;
        coeff[1520] <= 16'hb72d;
        coeff[1521] <= 16'hb765;
        coeff[1522] <= 16'hb79d;
        coeff[1523] <= 16'hb7d8;
        coeff[1524] <= 16'hb810;
        coeff[1525] <= 16'hb848;
        coeff[1526] <= 16'hb87d;
        coeff[1527] <= 16'hb8b5;
        coeff[1528] <= 16'hb8ed;
        coeff[1529] <= 16'hb922;
        coeff[1530] <= 16'hb95a;
        coeff[1531] <= 16'hb98e;
        coeff[1532] <= 16'hb9c3;
        coeff[1533] <= 16'hb9f8;
        coeff[1534] <= 16'hba2c;
        coeff[1535] <= 16'hba61;
        coeff[1536] <= 16'hba96;
        coeff[1537] <= 16'hbac7;
        coeff[1538] <= 16'hbafc;
        coeff[1539] <= 16'hbb2d;
        coeff[1540] <= 16'hbb5f;
        coeff[1541] <= 16'hbb90;
        coeff[1542] <= 16'hbbc5;
        coeff[1543] <= 16'hbbf6;
        coeff[1544] <= 16'hbc24;
        coeff[1545] <= 16'hbc56;
        coeff[1546] <= 16'hbc87;
        coeff[1547] <= 16'hbcb9;
        coeff[1548] <= 16'hbce7;
        coeff[1549] <= 16'hbd18;
        coeff[1550] <= 16'hbd46;
        coeff[1551] <= 16'hbd74;
        coeff[1552] <= 16'hbda6;
        coeff[1553] <= 16'hbdd4;
        coeff[1554] <= 16'hbe02;
        coeff[1555] <= 16'hbe30;
        coeff[1556] <= 16'hbe5e;
        coeff[1557] <= 16'hbe89;
        coeff[1558] <= 16'hbeb7;
        coeff[1559] <= 16'hbee5;
        coeff[1560] <= 16'hbf10;
        coeff[1561] <= 16'hbf3e;
        coeff[1562] <= 16'hbf69;
        coeff[1563] <= 16'hbf97;
        coeff[1564] <= 16'hbfc2;
        coeff[1565] <= 16'hbfed;
        coeff[1566] <= 16'hc018;
        coeff[1567] <= 16'hc043;
        coeff[1568] <= 16'hc06d;
        coeff[1569] <= 16'hc098;
        coeff[1570] <= 16'hc0c3;
        coeff[1571] <= 16'hc0ee;
        coeff[1572] <= 16'hc115;
        coeff[1573] <= 16'hc140;
        coeff[1574] <= 16'hc16b;
        coeff[1575] <= 16'hc193;
        coeff[1576] <= 16'hc1bd;
        coeff[1577] <= 16'hc1e5;
        coeff[1578] <= 16'hc20d;
        coeff[1579] <= 16'hc234;
        coeff[1580] <= 16'hc25f;
        coeff[1581] <= 16'hc286;
        coeff[1582] <= 16'hc2ae;
        coeff[1583] <= 16'hc2d5;
        coeff[1584] <= 16'hc2fd;
        coeff[1585] <= 16'hc325;
        coeff[1586] <= 16'hc34c;
        coeff[1587] <= 16'hc370;
        coeff[1588] <= 16'hc398;
        coeff[1589] <= 16'hc3bf;
        coeff[1590] <= 16'hc3e4;
        coeff[1591] <= 16'hc40b;
        coeff[1592] <= 16'hc42f;
        coeff[1593] <= 16'hc457;
        coeff[1594] <= 16'hc47b;
        coeff[1595] <= 16'hc4a3;
        coeff[1596] <= 16'hc4c7;
        coeff[1597] <= 16'hc4eb;
        coeff[1598] <= 16'hc513;
        coeff[1599] <= 16'hc537;
        coeff[1600] <= 16'hc55b;
        coeff[1601] <= 16'hc57f;
        coeff[1602] <= 16'hc5a4;
        coeff[1603] <= 16'hc5c8;
        coeff[1604] <= 16'hc5ec;
        coeff[1605] <= 16'hc610;
        coeff[1606] <= 16'hc635;
        coeff[1607] <= 16'hc659;
        coeff[1608] <= 16'hc67d;
        coeff[1609] <= 16'hc6a1;
        coeff[1610] <= 16'hc6c2;
        coeff[1611] <= 16'hc6e6;
        coeff[1612] <= 16'hc70b;
        coeff[1613] <= 16'hc72c;
        coeff[1614] <= 16'hc750;
        coeff[1615] <= 16'hc774;
        coeff[1616] <= 16'hc795;
        coeff[1617] <= 16'hc7b9;
        coeff[1618] <= 16'hc7da;
        coeff[1619] <= 16'hc7fe;
        coeff[1620] <= 16'hc81f;
        coeff[1621] <= 16'hc844;
        coeff[1622] <= 16'hc865;
        coeff[1623] <= 16'hc885;
        coeff[1624] <= 16'hc8aa;
        coeff[1625] <= 16'hc8cb;
        coeff[1626] <= 16'hc8ef;
        coeff[1627] <= 16'hc910;
        coeff[1628] <= 16'hc931;
        coeff[1629] <= 16'hc952;
        coeff[1630] <= 16'hc976;
        coeff[1631] <= 16'hc997;
        coeff[1632] <= 16'hc9b8;
        coeff[1633] <= 16'hc9d9;
        coeff[1634] <= 16'hc9fa;
        coeff[1635] <= 16'hca1e;
        coeff[1636] <= 16'hca3f;
        coeff[1637] <= 16'hca60;
        coeff[1638] <= 16'hca81;
        coeff[1639] <= 16'hcaa2;
        coeff[1640] <= 16'hcac3;
        coeff[1641] <= 16'hcae4;
        coeff[1642] <= 16'hcb05;
        coeff[1643] <= 16'hcb29;
        coeff[1644] <= 16'hcb4a;
        coeff[1645] <= 16'hcb6b;
        coeff[1646] <= 16'hcb8c;
        coeff[1647] <= 16'hcbad;
        coeff[1648] <= 16'hcbce;
        coeff[1649] <= 16'hcbee;
        coeff[1650] <= 16'hcc0f;
        coeff[1651] <= 16'hcc30;
        coeff[1652] <= 16'hcc51;
        coeff[1653] <= 16'hcc72;
        coeff[1654] <= 16'hcc93;
        coeff[1655] <= 16'hccb4;
        coeff[1656] <= 16'hccd8;
        coeff[1657] <= 16'hccf9;
        coeff[1658] <= 16'hcd1a;
        coeff[1659] <= 16'hcd3b;
        coeff[1660] <= 16'hcd5c;
        coeff[1661] <= 16'hcd7d;
        coeff[1662] <= 16'hcd9e;
        coeff[1663] <= 16'hcdbf;
        coeff[1664] <= 16'hcde3;
        coeff[1665] <= 16'hce04;
        coeff[1666] <= 16'hce25;
        coeff[1667] <= 16'hce46;
        coeff[1668] <= 16'hce67;
        coeff[1669] <= 16'hce88;
        coeff[1670] <= 16'hcea9;
        coeff[1671] <= 16'hceca;
        coeff[1672] <= 16'hceeb;
        coeff[1673] <= 16'hcf0c;
        coeff[1674] <= 16'hcf2d;
        coeff[1675] <= 16'hcf4e;
        coeff[1676] <= 16'hcf6e;
        coeff[1677] <= 16'hcf8f;
        coeff[1678] <= 16'hcfb0;
        coeff[1679] <= 16'hcfd1;
        coeff[1680] <= 16'hcff2;
        coeff[1681] <= 16'hd010;
        coeff[1682] <= 16'hd031;
        coeff[1683] <= 16'hd052;
        coeff[1684] <= 16'hd073;
        coeff[1685] <= 16'hd094;
        coeff[1686] <= 16'hd0b1;
        coeff[1687] <= 16'hd0d2;
        coeff[1688] <= 16'hd0f3;
        coeff[1689] <= 16'hd111;
        coeff[1690] <= 16'hd132;
        coeff[1691] <= 16'hd153;
        coeff[1692] <= 16'hd170;
        coeff[1693] <= 16'hd191;
        coeff[1694] <= 16'hd1af;
        coeff[1695] <= 16'hd1d0;
        coeff[1696] <= 16'hd1ee;
        coeff[1697] <= 16'hd20e;
        coeff[1698] <= 16'hd22c;
        coeff[1699] <= 16'hd24d;
        coeff[1700] <= 16'hd26b;
        coeff[1701] <= 16'hd28c;
        coeff[1702] <= 16'hd2a9;
        coeff[1703] <= 16'hd2c7;
        coeff[1704] <= 16'hd2e8;
        coeff[1705] <= 16'hd306;
        coeff[1706] <= 16'hd323;
        coeff[1707] <= 16'hd341;
        coeff[1708] <= 16'hd362;
        coeff[1709] <= 16'hd37f;
        coeff[1710] <= 16'hd39d;
        coeff[1711] <= 16'hd3bb;
        coeff[1712] <= 16'hd3d8;
        coeff[1713] <= 16'hd3f6;
        coeff[1714] <= 16'hd414;
        coeff[1715] <= 16'hd431;
        coeff[1716] <= 16'hd452;
        coeff[1717] <= 16'hd470;
        coeff[1718] <= 16'hd48a;
        coeff[1719] <= 16'hd4a8;
        coeff[1720] <= 16'hd4c6;
        coeff[1721] <= 16'hd4e3;
        coeff[1722] <= 16'hd501;
        coeff[1723] <= 16'hd51f;
        coeff[1724] <= 16'hd53c;
        coeff[1725] <= 16'hd55a;
        coeff[1726] <= 16'hd574;
        coeff[1727] <= 16'hd592;
        coeff[1728] <= 16'hd5af;
        coeff[1729] <= 16'hd5ca;
        coeff[1730] <= 16'hd5e7;
        coeff[1731] <= 16'hd605;
        coeff[1732] <= 16'hd61f;
        coeff[1733] <= 16'hd63d;
        coeff[1734] <= 16'hd657;
        coeff[1735] <= 16'hd675;
        coeff[1736] <= 16'hd68f;
        coeff[1737] <= 16'hd6ad;
        coeff[1738] <= 16'hd6c7;
        coeff[1739] <= 16'hd6e5;
        coeff[1740] <= 16'hd6ff;
        coeff[1741] <= 16'hd71a;
        coeff[1742] <= 16'hd737;
        coeff[1743] <= 16'hd752;
        coeff[1744] <= 16'hd76c;
        coeff[1745] <= 16'hd787;
        coeff[1746] <= 16'hd7a4;
        coeff[1747] <= 16'hd7bf;
        coeff[1748] <= 16'hd7d9;
        coeff[1749] <= 16'hd7f3;
        coeff[1750] <= 16'hd80e;
        coeff[1751] <= 16'hd828;
        coeff[1752] <= 16'hd842;
        coeff[1753] <= 16'hd85d;
        coeff[1754] <= 16'hd877;
        coeff[1755] <= 16'hd891;
        coeff[1756] <= 16'hd8ac;
        coeff[1757] <= 16'hd8c6;
        coeff[1758] <= 16'hd8dd;
        coeff[1759] <= 16'hd8f7;
        coeff[1760] <= 16'hd912;
        coeff[1761] <= 16'hd92c;
        coeff[1762] <= 16'hd943;
        coeff[1763] <= 16'hd95e;
        coeff[1764] <= 16'hd978;
        coeff[1765] <= 16'hd98f;
        coeff[1766] <= 16'hd9a9;
        coeff[1767] <= 16'hd9c0;
        coeff[1768] <= 16'hd9db;
        coeff[1769] <= 16'hd9f2;
        coeff[1770] <= 16'hda0c;
        coeff[1771] <= 16'hda23;
        coeff[1772] <= 16'hda3e;
        coeff[1773] <= 16'hda55;
        coeff[1774] <= 16'hda6c;
        coeff[1775] <= 16'hda83;
        coeff[1776] <= 16'hda9d;
        coeff[1777] <= 16'hdab4;
        coeff[1778] <= 16'hdacb;
        coeff[1779] <= 16'hdae2;
        coeff[1780] <= 16'hdaf9;
        coeff[1781] <= 16'hdb10;
        coeff[1782] <= 16'hdb27;
        coeff[1783] <= 16'hdb3f;
        coeff[1784] <= 16'hdb56;
        coeff[1785] <= 16'hdb6d;
        coeff[1786] <= 16'hdb84;
        coeff[1787] <= 16'hdb9b;
        coeff[1788] <= 16'hdbb2;
        coeff[1789] <= 16'hdbc6;
        coeff[1790] <= 16'hdbdd;
        coeff[1791] <= 16'hdbf4;
        coeff[1792] <= 16'hdc0b;
        coeff[1793] <= 16'hdc1f;
        coeff[1794] <= 16'hdc36;
        coeff[1795] <= 16'hdc49;
        coeff[1796] <= 16'hdc60;
        coeff[1797] <= 16'hdc74;
        coeff[1798] <= 16'hdc8b;
        coeff[1799] <= 16'hdc9f;
        coeff[1800] <= 16'hdcb3;
        coeff[1801] <= 16'hdcca;
        coeff[1802] <= 16'hdcde;
        coeff[1803] <= 16'hdcf1;
        coeff[1804] <= 16'hdd05;
        coeff[1805] <= 16'hdd19;
        coeff[1806] <= 16'hdd2d;
        coeff[1807] <= 16'hdd40;
        coeff[1808] <= 16'hdd54;
        coeff[1809] <= 16'hdd68;
        coeff[1810] <= 16'hdd7c;
        coeff[1811] <= 16'hdd90;
        coeff[1812] <= 16'hdda3;
        coeff[1813] <= 16'hddb7;
        coeff[1814] <= 16'hddcb;
        coeff[1815] <= 16'hdddb;
        coeff[1816] <= 16'hddef;
        coeff[1817] <= 16'hde03;
        coeff[1818] <= 16'hde13;
        coeff[1819] <= 16'hde27;
        coeff[1820] <= 16'hde3b;
        coeff[1821] <= 16'hde4b;
        coeff[1822] <= 16'hde5f;
        coeff[1823] <= 16'hde70;
        coeff[1824] <= 16'hde83;
        coeff[1825] <= 16'hde94;
        coeff[1826] <= 16'hdea4;
        coeff[1827] <= 16'hdeb8;
        coeff[1828] <= 16'hdec8;
        coeff[1829] <= 16'hded9;
        coeff[1830] <= 16'hdeed;
        coeff[1831] <= 16'hdefd;
        coeff[1832] <= 16'hdf0e;
        coeff[1833] <= 16'hdf1e;
        coeff[1834] <= 16'hdf2f;
        coeff[1835] <= 16'hdf3f;
        coeff[1836] <= 16'hdf50;
        coeff[1837] <= 16'hdf60;
        coeff[1838] <= 16'hdf70;
        coeff[1839] <= 16'hdf81;
        coeff[1840] <= 16'hdf91;
        coeff[1841] <= 16'hdfa2;
        coeff[1842] <= 16'hdfb2;
        coeff[1843] <= 16'hdfc3;
        coeff[1844] <= 16'hdfd3;
        coeff[1845] <= 16'hdfe0;
        coeff[1846] <= 16'hdff1;
        coeff[1847] <= 16'he001;
        coeff[1848] <= 16'he012;
        coeff[1849] <= 16'he01f;
        coeff[1850] <= 16'he030;
        coeff[1851] <= 16'he040;
        coeff[1852] <= 16'he04d;
        coeff[1853] <= 16'he05e;
        coeff[1854] <= 16'he06b;
        coeff[1855] <= 16'he07b;
        coeff[1856] <= 16'he088;
        coeff[1857] <= 16'he099;
        coeff[1858] <= 16'he0a6;
        coeff[1859] <= 16'he0b7;
        coeff[1860] <= 16'he0c4;
        coeff[1861] <= 16'he0d1;
        coeff[1862] <= 16'he0e1;
        coeff[1863] <= 16'he0ef;
        coeff[1864] <= 16'he0fc;
        coeff[1865] <= 16'he10c;
        coeff[1866] <= 16'he119;
        coeff[1867] <= 16'he127;
        coeff[1868] <= 16'he134;
        coeff[1869] <= 16'he144;
        coeff[1870] <= 16'he151;
        coeff[1871] <= 16'he15f;
        coeff[1872] <= 16'he16c;
        coeff[1873] <= 16'he179;
        coeff[1874] <= 16'he186;
        coeff[1875] <= 16'he197;
        coeff[1876] <= 16'he1a4;
        coeff[1877] <= 16'he1b1;
        coeff[1878] <= 16'he1be;
        coeff[1879] <= 16'he1cb;
        coeff[1880] <= 16'he1d8;
        coeff[1881] <= 16'he1e6;
        coeff[1882] <= 16'he1f3;
        coeff[1883] <= 16'he200;
        coeff[1884] <= 16'he20d;
        coeff[1885] <= 16'he217;
        coeff[1886] <= 16'he224;
        coeff[1887] <= 16'he231;
        coeff[1888] <= 16'he23f;
        coeff[1889] <= 16'he24c;
        coeff[1890] <= 16'he259;
        coeff[1891] <= 16'he266;
        coeff[1892] <= 16'he270;
        coeff[1893] <= 16'he27d;
        coeff[1894] <= 16'he28a;
        coeff[1895] <= 16'he298;
        coeff[1896] <= 16'he2a1;
        coeff[1897] <= 16'he2af;
        coeff[1898] <= 16'he2bc;
        coeff[1899] <= 16'he2c9;
        coeff[1900] <= 16'he2d3;
        coeff[1901] <= 16'he2e0;
        coeff[1902] <= 16'he2ed;
        coeff[1903] <= 16'he2f7;
        coeff[1904] <= 16'he304;
        coeff[1905] <= 16'he311;
        coeff[1906] <= 16'he31b;
        coeff[1907] <= 16'he328;
        coeff[1908] <= 16'he336;
        coeff[1909] <= 16'he340;
        coeff[1910] <= 16'he34d;
        coeff[1911] <= 16'he357;
        coeff[1912] <= 16'he364;
        coeff[1913] <= 16'he371;
        coeff[1914] <= 16'he37b;
        coeff[1915] <= 16'he388;
        coeff[1916] <= 16'he392;
        coeff[1917] <= 16'he39f;
        coeff[1918] <= 16'he3a9;
        coeff[1919] <= 16'he3b6;
        coeff[1920] <= 16'he3c3;
        coeff[1921] <= 16'he3cd;
        coeff[1922] <= 16'he3da;
        coeff[1923] <= 16'he3e4;
        coeff[1924] <= 16'he3ee;
        coeff[1925] <= 16'he3fb;
        coeff[1926] <= 16'he405;
        coeff[1927] <= 16'he412;
        coeff[1928] <= 16'he41c;
        coeff[1929] <= 16'he426;
        coeff[1930] <= 16'he430;
        coeff[1931] <= 16'he43d;
        coeff[1932] <= 16'he447;
        coeff[1933] <= 16'he451;
        coeff[1934] <= 16'he45b;
        coeff[1935] <= 16'he465;
        coeff[1936] <= 16'he472;
        coeff[1937] <= 16'he47c;
        coeff[1938] <= 16'he486;
        coeff[1939] <= 16'he490;
        coeff[1940] <= 16'he499;
        coeff[1941] <= 16'he4a3;
        coeff[1942] <= 16'he4ad;
        coeff[1943] <= 16'he4b7;
        coeff[1944] <= 16'he4c1;
        coeff[1945] <= 16'he4cb;
        coeff[1946] <= 16'he4d5;
        coeff[1947] <= 16'he4db;
        coeff[1948] <= 16'he4e5;
        coeff[1949] <= 16'he4ef;
        coeff[1950] <= 16'he4f9;
        coeff[1951] <= 16'he503;
        coeff[1952] <= 16'he50d;
        coeff[1953] <= 16'he513;
        coeff[1954] <= 16'he51d;
        coeff[1955] <= 16'he527;
        coeff[1956] <= 16'he52e;
        coeff[1957] <= 16'he538;
        coeff[1958] <= 16'he541;
        coeff[1959] <= 16'he548;
        coeff[1960] <= 16'he552;
        coeff[1961] <= 16'he55c;
        coeff[1962] <= 16'he562;
        coeff[1963] <= 16'he56c;
        coeff[1964] <= 16'he573;
        coeff[1965] <= 16'he57d;
        coeff[1966] <= 16'he583;
        coeff[1967] <= 16'he58d;
        coeff[1968] <= 16'he594;
        coeff[1969] <= 16'he59e;
        coeff[1970] <= 16'he5a4;
        coeff[1971] <= 16'he5ab;
        coeff[1972] <= 16'he5b5;
        coeff[1973] <= 16'he5bb;
        coeff[1974] <= 16'he5c5;
        coeff[1975] <= 16'he5cc;
        coeff[1976] <= 16'he5d2;
        coeff[1977] <= 16'he5dc;
        coeff[1978] <= 16'he5e3;
        coeff[1979] <= 16'he5e9;
        coeff[1980] <= 16'he5f0;
        coeff[1981] <= 16'he5fa;
        coeff[1982] <= 16'he601;
        coeff[1983] <= 16'he607;
        coeff[1984] <= 16'he60e;
        coeff[1985] <= 16'he618;
        coeff[1986] <= 16'he61e;
        coeff[1987] <= 16'he625;
        coeff[1988] <= 16'he62b;
        coeff[1989] <= 16'he632;
        coeff[1990] <= 16'he639;
        coeff[1991] <= 16'he642;
        coeff[1992] <= 16'he649;
        coeff[1993] <= 16'he650;
        coeff[1994] <= 16'he656;
        coeff[1995] <= 16'he65d;
        coeff[1996] <= 16'he663;
        coeff[1997] <= 16'he66a;
        coeff[1998] <= 16'he671;
        coeff[1999] <= 16'he677;
        coeff[2000] <= 16'he67e;
        coeff[2001] <= 16'he684;
        coeff[2002] <= 16'he68b;
        coeff[2003] <= 16'he691;
        coeff[2004] <= 16'he698;
        coeff[2005] <= 16'he69f;
        coeff[2006] <= 16'he6a5;
        coeff[2007] <= 16'he6ac;
        coeff[2008] <= 16'he6b2;
        coeff[2009] <= 16'he6b9;
        coeff[2010] <= 16'he6c0;
        coeff[2011] <= 16'he6c6;
        coeff[2012] <= 16'he6cd;
        coeff[2013] <= 16'he6d3;
        coeff[2014] <= 16'he6da;
        coeff[2015] <= 16'he6dd;
        coeff[2016] <= 16'he6e4;
        coeff[2017] <= 16'he6ea;
        coeff[2018] <= 16'he6f1;
        coeff[2019] <= 16'he6f8;
        coeff[2020] <= 16'he6fe;
        coeff[2021] <= 16'he705;
        coeff[2022] <= 16'he708;
        coeff[2023] <= 16'he70f;
        coeff[2024] <= 16'he715;
        coeff[2025] <= 16'he71c;
        coeff[2026] <= 16'he722;
        coeff[2027] <= 16'he729;
        coeff[2028] <= 16'he72c;
        coeff[2029] <= 16'he733;
        coeff[2030] <= 16'he739;
        coeff[2031] <= 16'he740;
        coeff[2032] <= 16'he747;
        coeff[2033] <= 16'he74d;
        coeff[2034] <= 16'he751;
        coeff[2035] <= 16'he757;
        coeff[2036] <= 16'he75e;
        coeff[2037] <= 16'he764;
        coeff[2038] <= 16'he768;
        coeff[2039] <= 16'he76e;
        coeff[2040] <= 16'he775;
        coeff[2041] <= 16'he77b;
        coeff[2042] <= 16'he782;
        coeff[2043] <= 16'he785;
        coeff[2044] <= 16'he78c;
        coeff[2045] <= 16'he792;
        coeff[2046] <= 16'he799;
        coeff[2047] <= 16'he7a0;
     end

   always @(posedge clk)
     val <= coeff[addr];

endmodule
